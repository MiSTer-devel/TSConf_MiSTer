-------------------------------------------------------------------[03.08.2014]
-- SDRAM Controller
-------------------------------------------------------------------------------
-- V1.0		03.08.2014	Initial release
-- modified for 8Mb SDRAM 15.03.2015 (Ivan Gorodetsky)

-- CLK		= 84 MHz	= 11.9 ns
-- WR/RD	= 5T		= 59.5 ns  
-- RFSH		= 6T		= 71.4 ns

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdram is
port(
	CLK		: in  std_logic;
	clk_28MHz: in  std_logic;
	c0 		: in  std_logic;
	c3 		: in  std_logic;

	-- Memory port
	loader	: in  std_logic;
	bsel  	: in  std_logic_vector(1  downto 0); -- Active HI
	A			: in  std_logic_vector(23 downto 0);
	DI			: in  std_logic_vector(15 downto 0);
	DO			: out std_logic_vector(15 downto 0);
	curr_cpu	: in  std_logic;
	DO_cpu	: out std_logic_vector(15 downto 0);
	REQ	 	: in  std_logic;
	RNW		: in  std_logic;

	-- SDRAM Pin
	CKE		: out std_logic;
	RAS_n		: out std_logic;
	CAS_n		: out std_logic;
	WE_n		: out std_logic;
	CS_n		: out std_logic;
	BA			: out std_logic_vector(1  downto 0);
	MA			: out std_logic_vector(12 downto 0);
	DQ			: inout std_logic_vector(15 downto 0);
	DQML		: out std_logic;
	DQMH		: out std_logic
);
end sdram;

architecture rtl of sdram is
	signal state 		: unsigned(4 downto 0) := "00000";
	signal col 			: std_logic_vector(7 downto 0);

	signal WR_in		: std_logic;
	signal RD_in		: std_logic;
	signal REQ_in		: std_logic;
	signal RNW_in		: std_logic;
	signal rd_op		: std_logic;
	signal RFSH_in		: std_logic;
	signal sdr_cmd		: std_logic_vector(2 downto 0);

	constant SdrCmd_xx 	: std_logic_vector(2 downto 0) := "111"; -- no operation
	constant SdrCmd_ac 	: std_logic_vector(2 downto 0) := "011"; -- activate
	constant SdrCmd_rd 	: std_logic_vector(2 downto 0) := "101"; -- read
	constant SdrCmd_wr 	: std_logic_vector(2 downto 0) := "100"; -- write		
	constant SdrCmd_pr 	: std_logic_vector(2 downto 0) := "010"; -- precharge all
	constant SdrCmd_re 	: std_logic_vector(2 downto 0) := "001"; -- refresh
	constant SdrCmd_ms 	: std_logic_vector(2 downto 0) := "000"; -- mode regiser set

-- Init-------------------------------------------------------------------		Idle		Read-------		Write------		Refresh-------
-- 00 01 02 03 04 05 06 07 08 09 0A 0B 0C 0D 0E 0F 10 11 12	13 14 15 16	17		18			19 1A 16 17		1B 1C 16 17		13 14 15 16 17
-- pr xx xx re xx xx xx xx xx xx re xx xx xx xx xx xx ms xx xx xx xx xx	xx		xx/ac/re	xx rd xx xx		xx wr xx xx		xx xx xx xx xx

begin

	process (clk_28MHz)
	begin 
		if rising_edge (clk_28MHz) then
			if c3 = '1' then --next_cycle
				RD_in		<= REQ and RNW;
				WR_in		<= REQ and not RNW;
				RFSH_in	<= not REQ;
			end if;

			if c0 = '1' then --NOT WORK
				RD_in 	<= '0';
				WR_in 	<= '0';
				RFSH_in 	<= '0';
			end if;
		end if;
	end process;
	
	process (CLK)
	begin
		if rising_edge(CLK) then
			---------------------------------------------------------				
			case state is
				-- Init
				when "00000" =>					-- s00
					sdr_cmd <= SdrCmd_pr;		-- PRECHARGE
					DQ <= (others => 'Z');
					MA <= (others => '1');
					BA <= "00";
					DQML <= '1';
					DQMH <= '1';
					state <= state + 1;

				when "00011" | "01010" =>		-- s03 s0A
					sdr_cmd <= SdrCmd_re;		-- REFRESH
					state <= state + 1;

				when "10001" =>					-- s11
					sdr_cmd <= SdrCmd_ms;		-- LOAD MODE REGISTER
					MA <= "000" & "1" & "00" & "010" & "0" & "000";				
					state <= state + 1;

				-- Idle		
				when "11000" =>					-- s18				
					rd_op <= '0';
					if rd_op = '1' then
						DO <= DQ;
						if curr_cpu = '1' then
							DO_cpu <= DQ;
						end if;
					end if;
					if RD_in = '1' or (WR_in = '1' and (loader = '1' or A(23) = '0')) then
						col <= A(7 downto 0);	-- LOCK COL
						sdr_cmd <= SdrCmd_ac;	-- ACTIVE
						BA <= A(10 downto 9);	
						MA <= "0"&A(23)&A(20 downto 11)&A(8);	-- RAW_ADDR(12..0)
						DQML <= not (bsel(0) or RD_in);
						DQMH <= not (bsel(1) or RD_in);
						rd_op <= RD_in;
						state <= state + 1;
					elsif RFSH_in = '1' then
						sdr_cmd <= SdrCmd_re;	-- REFRESH
						state <= "10011";			-- s13
					end if;

				-- A24 A23 A22 A21 A20 A19 A18 A17 A16 A15 A14 A13 A12 A11 A10 A9 A8 A7 A6 A5 A4 A3 A2 A1 A0
				-- -----------------------ROW------------------------- BA1 BA0 -----------COLUMN------------		

				-- Single read/write - with auto precharge
				when "11010" =>					-- s1A
					MA <= "00100" & col; 		-- A10 = 1 enable auto precharge; A9..0 = column
					state <= "10110";				-- s16
					if rd_op = '1' then
						sdr_cmd <= SdrCmd_rd;	-- READ
					else
						sdr_cmd <= SdrCmd_wr;	-- WRITE
						DQ <= DI;
					end if;
					
				when others =>
					DQ <= (others => 'Z');
					sdr_cmd <= SdrCmd_xx;		-- NOP
					state <= state + 1;
			end case;
		end if;
	end process;

	CKE 	<= '1';
	CS_n  <= '0';
	RAS_n <= sdr_cmd(2);
	CAS_n <= sdr_cmd(1);
	WE_n 	<= sdr_cmd(0);

end rtl;